`timescale 1ns / 1ps
module StallControlLogic(
    input [31:0]inst_in,
    input [31:0]Data_in,

    output id_shouldStall
    );
    
endmodule